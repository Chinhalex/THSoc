
module system (
	clk_clk,
	red_leds_0_conduit_end_export,
	reset_reset_n,
	switches_0_conduit_end_export);	

	input		clk_clk;
	output	[31:0]	red_leds_0_conduit_end_export;
	input		reset_reset_n;
	input	[31:0]	switches_0_conduit_end_export;
endmodule
