// system_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system_tb (
	);

	wire         system_inst_clk_bfm_clk_clk;                           // system_inst_clk_bfm:clk -> [system_inst:clk_clk, system_inst_red_leds_0_conduit_end_bfm:clk, system_inst_reset_bfm:clk, system_inst_switches_0_conduit_end_bfm:clk]
	wire  [31:0] system_inst_red_leds_0_conduit_end_export;             // system_inst:red_leds_0_conduit_end_export -> system_inst_red_leds_0_conduit_end_bfm:sig_export
	wire  [31:0] system_inst_switches_0_conduit_end_bfm_conduit_export; // system_inst_switches_0_conduit_end_bfm:sig_export -> system_inst:switches_0_conduit_end_export
	wire         system_inst_reset_bfm_reset_reset;                     // system_inst_reset_bfm:reset -> [system_inst:reset_reset_n, system_inst_red_leds_0_conduit_end_bfm:reset, system_inst_switches_0_conduit_end_bfm:reset]

	system system_inst (
		.clk_clk                       (system_inst_clk_bfm_clk_clk),                           //                    clk.clk
		.red_leds_0_conduit_end_export (system_inst_red_leds_0_conduit_end_export),             // red_leds_0_conduit_end.export
		.reset_reset_n                 (system_inst_reset_bfm_reset_reset),                     //                  reset.reset_n
		.switches_0_conduit_end_export (system_inst_switches_0_conduit_end_bfm_conduit_export)  // switches_0_conduit_end.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) system_inst_clk_bfm (
		.clk (system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm system_inst_red_leds_0_conduit_end_bfm (
		.clk        (system_inst_clk_bfm_clk_clk),               //     clk.clk
		.reset      (~system_inst_reset_bfm_reset_reset),        //   reset.reset
		.sig_export (system_inst_red_leds_0_conduit_end_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) system_inst_reset_bfm (
		.reset (system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 system_inst_switches_0_conduit_end_bfm (
		.clk        (system_inst_clk_bfm_clk_clk),                           //     clk.clk
		.reset      (~system_inst_reset_bfm_reset_reset),                    //   reset.reset
		.sig_export (system_inst_switches_0_conduit_end_bfm_conduit_export)  // conduit.export
	);

endmodule
